

module portevent(
);


endmodule