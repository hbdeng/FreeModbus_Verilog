

module portserial(
    // inputs
    inMBPortSerialEnable,
    inMBPortSerialInit,
    inMBPortSerialPutByte,
    inMBPortSerialGetByte,
    inRxEnable,
    inTxEnable,
    
    // inouts
    
    // outpus
    outUARTTxReadyISR,
    outUARTRxISR
);

    /**
     * Put uart module here
     **/

endmodule