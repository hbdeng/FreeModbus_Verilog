module demo(

);

endmodule