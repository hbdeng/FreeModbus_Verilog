

module porttimer(
    // inputs
    inMBPortTimersInit,
    inMBPortTimersEnable,
    inMBPortTimersDisable,
    
    // inouts
    
    // outpus
    outTIMERExpiredISR
);


endmodule
